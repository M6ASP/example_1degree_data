netcdf ocean.static {
dimensions:
	yq = 320 ;
	xq = 360 ;
	yh = 320 ;
	xh = 360 ;
variables:
	float Coriolis(yq, xq) ;
		Coriolis:long_name = "Coriolis parameter at corner (Bu) points" ;
		Coriolis:units = "s-1" ;
		Coriolis:missing_value = 1.e+20f ;
		Coriolis:_FillValue = 1.e+20f ;
		Coriolis:cell_methods = "time: point" ;
		Coriolis:interp_method = "none" ;
	float area_t(yh, xh) ;
		area_t:long_name = "Surface area of tracer (T) cells" ;
		area_t:units = "m2" ;
		area_t:missing_value = 1.e+20f ;
		area_t:_FillValue = 1.e+20f ;
		area_t:cell_methods = "area:sum yh:sum xh:sum time: point" ;
	float areacello(yh, xh) ;
		areacello:long_name = "Ocean Grid-Cell Area" ;
		areacello:units = "m2" ;
		areacello:missing_value = 1.e+20f ;
		areacello:_FillValue = 1.e+20f ;
		areacello:cell_methods = "area:sum yh:sum xh:sum time: point" ;
		areacello:standard_name = "cell_area" ;
	float areacello_bu(yq, xq) ;
		areacello_bu:long_name = "Ocean Grid-Cell Area" ;
		areacello_bu:units = "m2" ;
		areacello_bu:missing_value = 1.e+20f ;
		areacello_bu:_FillValue = 1.e+20f ;
		areacello_bu:cell_methods = "area:sum yq:sum xq:sum time: point" ;
		areacello_bu:standard_name = "cell_area" ;
	float areacello_cu(yh, xq) ;
		areacello_cu:long_name = "Ocean Grid-Cell Area" ;
		areacello_cu:units = "m2" ;
		areacello_cu:missing_value = 1.e+20f ;
		areacello_cu:_FillValue = 1.e+20f ;
		areacello_cu:cell_methods = "area:sum yh:sum xq:sum time: point" ;
		areacello_cu:standard_name = "cell_area" ;
	float areacello_cv(yq, xh) ;
		areacello_cv:long_name = "Ocean Grid-Cell Area" ;
		areacello_cv:units = "m2" ;
		areacello_cv:missing_value = 1.e+20f ;
		areacello_cv:_FillValue = 1.e+20f ;
		areacello_cv:cell_methods = "area:sum yq:sum xh:sum time: point" ;
		areacello_cv:standard_name = "cell_area" ;
	float depth_ocean(yh, xh) ;
		depth_ocean:long_name = "Depth of the ocean at tracer points" ;
		depth_ocean:units = "m" ;
		depth_ocean:missing_value = 1.e+20f ;
		depth_ocean:_FillValue = 1.e+20f ;
		depth_ocean:cell_methods = "area:mean yh:mean xh:mean time: point" ;
		depth_ocean:cell_measures = "area: area_t" ;
		depth_ocean:standard_name = "sea_floor_depth_below_geoid" ;
	float deptho(yh, xh) ;
		deptho:long_name = "Sea Floor Depth" ;
		deptho:units = "m" ;
		deptho:missing_value = 1.e+20f ;
		deptho:_FillValue = 1.e+20f ;
		deptho:cell_methods = "area:mean yh:mean xh:mean time: point" ;
		deptho:cell_measures = "area: area_t" ;
		deptho:standard_name = "sea_floor_depth_below_geoid" ;
	float dxCu(yh, xq) ;
		dxCu:long_name = "Delta(x) at u points (meter)" ;
		dxCu:units = "m" ;
		dxCu:missing_value = 1.e+20f ;
		dxCu:_FillValue = 1.e+20f ;
		dxCu:cell_methods = "time: point" ;
		dxCu:interp_method = "none" ;
	float dxCv(yq, xh) ;
		dxCv:long_name = "Delta(x) at v points (meter)" ;
		dxCv:units = "m" ;
		dxCv:missing_value = 1.e+20f ;
		dxCv:_FillValue = 1.e+20f ;
		dxCv:cell_methods = "time: point" ;
		dxCv:interp_method = "none" ;
	float dxt(yh, xh) ;
		dxt:long_name = "Delta(x) at thickness/tracer points (meter)" ;
		dxt:units = "m" ;
		dxt:missing_value = 1.e+20f ;
		dxt:_FillValue = 1.e+20f ;
		dxt:cell_methods = "time: point" ;
		dxt:interp_method = "none" ;
	float dyCu(yh, xq) ;
		dyCu:long_name = "Delta(y) at u points (meter)" ;
		dyCu:units = "m" ;
		dyCu:missing_value = 1.e+20f ;
		dyCu:_FillValue = 1.e+20f ;
		dyCu:cell_methods = "time: point" ;
		dyCu:interp_method = "none" ;
	float dyCv(yq, xh) ;
		dyCv:long_name = "Delta(y) at v points (meter)" ;
		dyCv:units = "m" ;
		dyCv:missing_value = 1.e+20f ;
		dyCv:_FillValue = 1.e+20f ;
		dyCv:cell_methods = "time: point" ;
		dyCv:interp_method = "none" ;
	float dyt(yh, xh) ;
		dyt:long_name = "Delta(y) at thickness/tracer points (meter)" ;
		dyt:units = "m" ;
		dyt:missing_value = 1.e+20f ;
		dyt:_FillValue = 1.e+20f ;
		dyt:cell_methods = "time: point" ;
		dyt:interp_method = "none" ;
	float geolat(yh, xh) ;
		geolat:long_name = "Latitude of tracer (T) points" ;
		geolat:units = "degrees_north" ;
		geolat:missing_value = 1.e+20f ;
		geolat:_FillValue = 1.e+20f ;
		geolat:cell_methods = "time: point" ;
	float geolat_c(yq, xq) ;
		geolat_c:long_name = "Latitude of corner (Bu) points" ;
		geolat_c:units = "degrees_north" ;
		geolat_c:missing_value = 1.e+20f ;
		geolat_c:_FillValue = 1.e+20f ;
		geolat_c:cell_methods = "time: point" ;
		geolat_c:interp_method = "none" ;
	float geolat_u(yh, xq) ;
		geolat_u:long_name = "Latitude of zonal velocity (Cu) points" ;
		geolat_u:units = "degrees_north" ;
		geolat_u:missing_value = 1.e+20f ;
		geolat_u:_FillValue = 1.e+20f ;
		geolat_u:cell_methods = "time: point" ;
		geolat_u:interp_method = "none" ;
	float geolat_v(yq, xh) ;
		geolat_v:long_name = "Latitude of meridional velocity (Cv) points" ;
		geolat_v:units = "degrees_north" ;
		geolat_v:missing_value = 1.e+20f ;
		geolat_v:_FillValue = 1.e+20f ;
		geolat_v:cell_methods = "time: point" ;
		geolat_v:interp_method = "none" ;
	float geolon(yh, xh) ;
		geolon:long_name = "Longitude of tracer (T) points" ;
		geolon:units = "degrees_east" ;
		geolon:missing_value = 1.e+20f ;
		geolon:_FillValue = 1.e+20f ;
		geolon:cell_methods = "time: point" ;
	float geolon_c(yq, xq) ;
		geolon_c:long_name = "Longitude of corner (Bu) points" ;
		geolon_c:units = "degrees_east" ;
		geolon_c:missing_value = 1.e+20f ;
		geolon_c:_FillValue = 1.e+20f ;
		geolon_c:cell_methods = "time: point" ;
		geolon_c:interp_method = "none" ;
	float geolon_u(yh, xq) ;
		geolon_u:long_name = "Longitude of zonal velocity (Cu) points" ;
		geolon_u:units = "degrees_east" ;
		geolon_u:missing_value = 1.e+20f ;
		geolon_u:_FillValue = 1.e+20f ;
		geolon_u:cell_methods = "time: point" ;
		geolon_u:interp_method = "none" ;
	float geolon_v(yq, xh) ;
		geolon_v:long_name = "Longitude of meridional velocity (Cv) points" ;
		geolon_v:units = "degrees_east" ;
		geolon_v:missing_value = 1.e+20f ;
		geolon_v:_FillValue = 1.e+20f ;
		geolon_v:cell_methods = "time: point" ;
		geolon_v:interp_method = "none" ;
	float sftof(yh, xh) ;
		sftof:long_name = "Sea Area Fraction" ;
		sftof:units = "%" ;
		sftof:missing_value = 1.e+20f ;
		sftof:_FillValue = 1.e+20f ;
		sftof:cell_methods = "area:mean yh:mean xh:mean time: point" ;
		sftof:standard_name = "SeaAreaFraction" ;
	float wet(yh, xh) ;
		wet:long_name = "0 if land, 1 if ocean at tracer points" ;
		wet:units = "none" ;
		wet:missing_value = 1.e+20f ;
		wet:_FillValue = 1.e+20f ;
		wet:cell_methods = "time: point" ;
		wet:cell_measures = "area: area_t" ;
	float wet_c(yq, xq) ;
		wet_c:long_name = "0 if land, 1 if ocean at corner (Bu) points" ;
		wet_c:units = "none" ;
		wet_c:missing_value = 1.e+20f ;
		wet_c:_FillValue = 1.e+20f ;
		wet_c:cell_methods = "time: point" ;
		wet_c:interp_method = "none" ;
	float wet_u(yh, xq) ;
		wet_u:long_name = "0 if land, 1 if ocean at zonal velocity (Cu) points" ;
		wet_u:units = "none" ;
		wet_u:missing_value = 1.e+20f ;
		wet_u:_FillValue = 1.e+20f ;
		wet_u:cell_methods = "time: point" ;
		wet_u:interp_method = "none" ;
	float wet_v(yq, xh) ;
		wet_v:long_name = "0 if land, 1 if ocean at meridional velocity (Cv) points" ;
		wet_v:units = "none" ;
		wet_v:missing_value = 1.e+20f ;
		wet_v:_FillValue = 1.e+20f ;
		wet_v:cell_methods = "time: point" ;
		wet_v:interp_method = "none" ;
	double xh(xh) ;
		xh:long_name = "h point nominal longitude" ;
		xh:units = "degrees_east" ;
		xh:cartesian_axis = "X" ;
	double xq(xq) ;
		xq:long_name = "q point nominal longitude" ;
		xq:units = "degrees_east" ;
		xq:cartesian_axis = "X" ;
	double yh(yh) ;
		yh:long_name = "h point nominal latitude" ;
		yh:units = "degrees_north" ;
		yh:cartesian_axis = "Y" ;
	double yq(yq) ;
		yq:long_name = "q point nominal latitude" ;
		yq:units = "degrees_north" ;
		yq:cartesian_axis = "Y" ;

// global attributes:
		:filename = "ocean.static.nc" ;
		:title = "SPEAR_c96_o1_Control_1850_E50" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:external_variables = "area_t area_t area_t" ;
}
